module instruction_Mem (
        input   [31:0] address
    ,   input   [31:0] instr_in
    ,   output  [31:0] instr_ID
    ,   output         start
);
    
endmodule
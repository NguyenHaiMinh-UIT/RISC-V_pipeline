module loadhazard (
    input [4:0] rs1D,
    input [4:0] rs2D,
    input [4:0] rdE,
    input [1:0] write_back_E,
    output stallF,
    output stallD,
    output FlushE
);
    
endmodule
module harzard_unit (
        input rs1
    ,   input rs2
    ,   input rdE
    ,   output Stall_ID
    ,   output Stall_IF
    ,   output Flush_IE
    ,   output WriteBack_EX
);
    
endmodule
module harzard_unit (
    input in,
    output out
);
    
endmodule
module pc (
        input clk,rst
    ,   input   [31:0]  pcF
    ,   output  [31:0]  pc_plus4
);
    
endmodule
module signExtend (
        input   [31:7]  instr_D
    ,   input           immD
    ,   output  [31:0]  imm_out_D
);
    
endmodule